module clock_divisor_nopara(clk1, clk);
input clk;
output clk1;
reg [1:0] num;
wire [1:0] next_num;

always @(posedge clk) begin
  num <= next_num;
end

assign next_num = num + 1'b1;
assign clk1 = num[1];
endmodule
